
interface ahb_interface(input clk, input rst_n);

   logic [31:0]  addr;

endinterface
